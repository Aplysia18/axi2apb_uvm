`ifndef RESET_PKG_SV
`define RESET_PKG_SV

`include "../public/reset_vip/reset_tr.sv"
`include "../public/reset_vip/reset_vif.sv"
`include "../public/reset_vip/reset_agent.sv"

`endif  // AXI_PKG_SV
